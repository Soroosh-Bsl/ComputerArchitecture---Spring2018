module rom(address,data, reset);
input [9:0] address; //needs to be changed
input reset;
output [25:0] data;	//needs to be changed
reg [25:0] array[300:0];	//needs to be changed

// 1234567890
always @(negedge reset)
begin
//fetch = 0
array[0] = 26'b00001_00001_000_000_0000000000;//PC to AR, INCPC
array[1] = 26'b00010_00000_000_000_0000000000;//READ MEM
array[2] = 26'b01111_00000_000_000_0000000000;//loadIR
array[3] = 26'b00000_00000_111_000_0000000000;//GOTO MAP

//iadd = 4
array[4] = 26'b00011_00010_000_000_0000000000;//SP_STAR to AR, decSP
array[5] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[6] = 26'b00000_01100_000_000_0000000000;//loadOP
array[7] = 26'b00011_00010_000_000_0000000000;//SP_STAR to AR, decSP
array[8] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[9] = 26'b00100_00000_000_000_0000000000;//loadDR
array[10] = 26'b11000_00011_000_000_0000000000;//SP to AR, RES+
array[11] = 26'b00101_00000_000_000_0000000000;//RES to mem
array[12] = 26'b00000_00100_110_000_0000000000;//incSP

//isub = 13
array[10+3] = 26'b00011_00010_000_000_0000000000;//SP_STAR to AR, decSP
array[10+4] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[10+5] = 26'b00000_01100_000_000_0000000000;//loadOP
array[10+6] = 26'b00011_00010_000_000_0000000000;//SP_STAR to AR, decSP
array[10+7] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[10+8] = 26'b00100_00000_000_000_0000000000;//loadDR
array[10+9] = 26'b11000_01111_000_000_0000000000;//SP to AR, RES-
array[10+10] = 26'b00101_00000_000_000_0000000000;//RES to mem
array[10+11] = 26'b00000_00100_110_000_0000000000;//incSP

//iand = 22
array[19+3] = 26'b00011_00010_000_000_0000000000;//SP_STAR to AR, decSP
array[19+4] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[19+5] = 26'b00000_01100_000_000_0000000000;//loadOP
array[19+6] = 26'b00011_00010_000_000_0000000000;//SP_STAR to AR, decSP
array[19+7] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[19+8] = 26'b00100_00000_000_000_0000000000;//loadDR
array[19+9] = 26'b11000_01010_000_000_0000000000;//SP to AR, RES MULT
array[19+10] = 26'b00101_00000_000_000_0000000000;//RES to mem
array[19+11] = 26'b00000_00100_110_000_0000000000;//incSP

//ior = 31
array[28+3] = 26'b00011_00010_000_000_0000000000;//SP_STAR to AR, decSP
array[28+4] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[28+5] = 26'b00000_01100_000_000_0000000000;//loadOP
array[28+6] = 26'b00011_00010_000_000_0000000000;//SP_STAR to AR, decSP
array[28+7] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[28+8] = 26'b00100_00000_000_000_0000000000;//loadDR
array[28+9] = 26'b11000_01011_000_000_0000000000;//SP to AR, RES OR
array[28+10] = 26'b00101_00000_000_000_0000000000;//RES to mem
array[28+11] = 26'b00000_00100_110_000_0000000000;//incSP

//GOTO = 40
array[37+3] = 26'b00001_00101_000_000_0000000000;//PC to AR, PC+TWO
array[37+4] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[37+5] = 26'b00100_00000_000_000_0000000000;//loadDR
array[37+6] = 26'b00000_00110_000_000_0000000000;//DR to PC branch

//IFEQ = 44
array[41+3] = 26'b00011_00010_000_000_0000000000;//SP_STAR to AR, decSP
array[41+4] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[41+5] = 26'b00100_00000_001_000_0000101111;//loadDR, if Z then to SEVEN %%%%%%%%%
array[41+6] = 26'b00000_00101_110_000_0000000000;//PC+TWO, FINISH to Fetch
array[41+7] = 26'b00001_00101_000_000_0000000000;//PC to AR, PC+TWO
array[41+8] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[41+9] = 26'b00000_00111_110_000_0000000000;//loadPC branch memory

//IFLT = 51
array[48+3] = 26'b00011_00010_000_000_0000000000;//SP_STAR to AR, decSP
array[48+4] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[48+5] = 26'b00100_00000_001_001_0000110110;//loadDR, if N then to SEVEN %%%%%%%%%
array[48+6] = 26'b00000_00101_110_000_0000000000;//PC+TWO, FINISH to Fetch
array[48+7] = 26'b00001_00101_000_000_0000000000;//PC to AR, PC+TWO
array[48+8] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[48+9] = 26'b00000_00111_110_000_0000000000;//loadPC branch memory

//IF_ICMPEQ = 58
array[55+3] = 26'b00011_00010_000_000_0000000000;//SP_STAR to AR, decSP
array[55+4] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[55+5] = 26'b00100_00000_000_000_0000000000;//loadDR
array[55+6] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[55+7] = 26'b00000_01100_000_000_0000000000;//loadOP
array[55+8] = 26'b00000_01111_001_000_0001000000;//RES-, if Z to TEN %%%%%%%%%%%
array[55+9] = 26'b00000_00101_110_000_0000000000;//PC+TWO, FINISH to Fetch
array[55+10] = 26'b00001_00101_000_000_0000000000;//PC to AR, PC+TWO
array[55+11] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[55+12] = 26'b00000_00111_110_000_0000000000;//loadPC branch memory

//NOP = 68
array[65+3] = 26'b00000_00000_110_000_0000000000;//

//POP = 69
array[66+3] = 26'b00000_00010_110_000_0000000000;//decSP

//dup = 70 OK
array[67+3] = 26'b00011_00000_000_000_0000000000;//SP_STAR to AR
array[67+4] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[67+5] = 26'b00100_00000_000_000_0000000000;//loadDR
array[67+6] = 26'b11000_00100_000_000_0000000000;//SP to AR, incSP
array[67+7] = 26'b00110_00000_110_000_0000000000;//DR to mem

//iload __TWO__ = 75
array[72+3] = 26'b00001_00101_000_000_0000000000;//PC to AR, PC+TWO
array[72+4] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[72+5] = 26'b00000_01100_000_000_0000000000;//loadOP
array[72+6] = 26'b00000_01001_000_000_0000000000;//OP<<TWO
array[72+7] = 26'b01001_00000_000_000_0000000000;//LV to DR
array[72+8] = 26'b00000_00011_000_000_0000000000;//RES+
array[72+9] = 26'b01010_00000_000_000_0000000000;//RES to AR
array[72+10] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[72+11] = 26'b00100_00000_000_000_0000000000;//loadDR
array[72+12] = 26'b11000_00100_000_000_0000000000;//SP to AR, incSP
array[72+13] = 26'b00110_00000_110_000_0000000000;//DR to mem

//iload __ONE__ = 86
array[83+3] = 26'b00001_00001_000_000_0000000000;//PC to AR, PC+ONE
array[83+4] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[83+5] = 26'b00000_01100_000_000_0000000000;//loadOP
array[83+6] = 26'b00000_01001_000_000_0000000000;//OP<<TWO
array[83+7] = 26'b01001_00000_000_000_0000000000;//LV to DR
array[83+8] = 26'b00000_00011_000_000_0000000000;//RES+
array[83+9] = 26'b01010_00000_000_000_0000000000;//RES to AR
array[83+10] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[83+11] = 26'b00100_00000_000_000_0000000000;//loadDR
array[83+12] = 26'b11000_00100_000_000_0000000000;//SP to AR, incSP
array[83+13] = 26'b00110_00000_110_000_0000000000;//DR to mem

//istore __TWO__ = 97
array[94+3] = 26'b00011_00010_000_000_0000000000;//SP_STAR to AR, decSP
array[94+4] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[94+5] = 26'b00111_00000_000_000_0000000000;//loadTR
array[94+6] = 26'b00001_00101_000_000_0000000000;//PC to AR, PC+TWO
array[94+7] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[94+8] = 26'b00000_01100_000_000_0000000000;//loadOP
array[94+9] = 26'b00000_01001_000_000_0000000000;//OP<<TWO
array[94+10] = 26'b01001_00000_000_000_0000000000;//LV to DR
array[94+11] = 26'b00000_00011_000_000_0000000000;//RES+
array[94+12] = 26'b01010_00000_000_000_0000000000;//RES to AR
array[94+13] = 26'b01000_00000_110_000_0000000000;//TR to mem

//istore __ONE__ = 108
array[105+3] = 26'b00011_00010_000_000_0000000000;//SP_STAR to AR, decSP
array[105+4] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[105+5] = 26'b00111_00000_000_000_0000000000;//loadTR
array[105+6] = 26'b00001_00101_000_000_0000000000;//PC to AR, PC+TWO
array[105+7] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[105+8] = 26'b00000_01100_000_000_0000000000;//loadOP
array[105+9] = 26'b00000_01001_000_000_0000000000;//OP<<TWO
array[105+10] = 26'b01001_00000_000_000_0000000000;//LV to DR
array[105+11] = 26'b00000_00011_000_000_0000000000;//RES+
array[105+12] = 26'b01010_00000_000_000_0000000000;//RES to AR
array[105+13] = 26'b01000_00000_110_000_0000000000;//TR to mem

//bipush __TWO__ = 119
array[116+3] = 26'b00001_00101_000_000_0000000000;//PC to AR, PC+TWO
array[116+4] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[116+5] = 26'b00100_00000_000_000_0000000000;//loadDR
array[116+6] = 26'b11000_00100_000_000_0000000000;//SP to AR, incSP
array[116+7] = 26'b00110_00000_110_000_0000000000;//DR to mem

//bipush __ONE__ = 130
array[127+3] = 26'b00001_00001_000_000_0000000000;//PC to AR, PC+ONE
array[127+4] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[127+5] = 26'b00100_00000_000_000_0000000000;//loadDR
array[127+6] = 26'b11000_00100_000_000_0000000000;//SP to AR, incSP
array[127+7] = 26'b00110_00000_110_000_0000000000;//DR to mem

//SWAP = 141
array[138+3] = 26'b00011_00010_000_000_0000000000;//SP_STAR to AR, decSP
array[138+4] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[138+5] = 26'b00000_01100_000_000_0000000000;//loadOP
array[138+6] = 26'b00011_00010_000_000_0000000000;//SP_STAR to AR, decSP
array[138+7] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[138+8] = 26'b00100_00000_000_000_0000000000;//loadDR
array[138+9] = 26'b11000_00100_000_000_0000000000;//SP to AR, incSP
array[138+10] = 26'b00000_10000_000_000_0000000000;//OP to RESULT
array[138+11] = 26'b00101_00000_000_000_0000000000;//RES to mem
array[138+12] = 26'b11000_00100_000_000_0000000000;//SP to AR, incSP
array[138+13] = 26'b00110_00000_110_000_0000000000;//DR to mem

//wide = 152
array[149+3] = 26'b00000_00000_110_111_0000000000;

//ldc_w = 153
array[150+3] = 26'b00001_00101_000_000_0000000000;//PC to AR, PC+TWO
array[150+4] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[150+5] = 26'b00000_01100_000_000_0000000000;//loadOP
array[150+6] = 26'b00000_01001_000_000_0000000000;//OP<<TWO
array[150+7] = 26'b01110_00000__000_000_0000000000;//CPP to DR
array[150+8] = 26'b00000_00011_000_000_0000000000;//RES+
array[150+9] = 26'b01010_00000_000_000_0000000000;//RES to AR
array[150+10] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[150+11] = 26'b00000_01100_000_000_0000000000;//loadOP
array[150+12] = 26'b11000_00100_000_000_0000000000;//SP to AR, incSP
array[150+13] = 26'b00000_10000_000_000_0000000000;//OP to RESULT
array[150+14] = 26'b00101_00000_110_000_0000000000;//RES to mem

//inc = 165
array[162+3] = 26'b00001_00101_000_000_0000000000;//PC to AR, PC+TWO
array[162+4] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[162+5] = 26'b00000_01100_000_000_0000000000;//loadOP
array[162+6] = 26'b00000_01001_000_000_0000000000;//OP<<TWO
array[162+7] = 26'b01001_00000_000_000_0000000000;//LV to DR
array[162+8] = 26'b00000_00011_000_000_0000000000;//RES+
array[162+9] = 26'b01010_00000_000_000_0000000000;//RES to AR
array[162+10] = 26'b01011_00000_000_000_0000000000;//RES to TR
array[162+11] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[162+12] = 26'b00100_00000_000_000_0000000000;//loadDR
array[162+13] = 26'b00001_00001_000_000_0000000000;//PC to AR, PC+ONE
array[162+14] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[162+15] = 26'b00000_01100_000_000_0000000000;//loadOP
array[162+16] = 26'b00000_00011_000_000_0000000000;//RES+
array[162+17] = 26'b11100_00000_000_000_0000000000;//TR to AR
array[162+18] = 26'b00101_00000_110_000_0000000000;//RES to mem

//inc __TWO__= 240
array[237+3] = 26'b00001_00101_000_000_0000000000;//PC to AR, PC+TWO
array[237+4] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[237+5] = 26'b00000_01100_000_000_0000000000;//loadOP
array[237+6] = 26'b00000_01001_000_000_0000000000;//OP<<TWO
array[237+7] = 26'b01001_00000_000_000_0000000000;//LV to DR
array[237+8] = 26'b00000_00011_000_000_0000000000;//RES+
array[237+9] = 26'b01010_00000_000_000_0000000000;//RES to AR
array[237+10] = 26'b01011_00000_000_000_0000000000;//RES to TR
array[237+11] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[237+12] = 26'b00100_00000_000_000_0000000000;//loadDR
array[237+13] = 26'b00001_00101_000_000_0000000000;//PC to AR, PC+TWO
array[237+14] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[237+15] = 26'b00000_01100_000_000_0000000000;//loadOP
array[237+16] = 26'b00000_00011_000_000_0000000000;//RES+
array[237+17] = 26'b11100_00000_000_000_0000000000;//TR to AR
array[237+18] = 26'b00101_00000_110_000_0000000000;//RES to mem

//invoke = 181
array[178+3] = 26'b00001_00101_000_000_0000000000;//PC to AR, PC+TWO
array[178+4] = 26'b01100_00000_000_000_0000000000;//PC to SR
array[178+5] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[178+6] = 26'b00000_01100_000_000_0000000000;//loadOP
array[178+7] = 26'b00000_01001_000_000_0000000000;//OP<<TWO
array[178+8] = 26'b01110_00000__000_000_0000000000;//CPP to DR
array[178+9] = 26'b00000_00011_000_000_0000000000;//RES+
array[178+10] = 26'b01010_00000_000_000_0000000000;//RES to AR
array[178+11] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[178+12] = 26'b00000_11111_000_000_0000000000;//reloadPC from mem
array[178+13] = 26'b10011_00000_000_000_0000000000;//PC to TR

array[178+14] = 26'b00001_00101_000_000_0000000000;//PC to AR, PC+TWO
array[178+15] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[178+16] = 26'b00000_01100_000_000_0000000000;//loadOP
array[178+17] = 26'b00000_01001_000_000_0000000000;//OP<<TWO
array[178+18] = 26'b10001_00000_000_000_0000000000;//SP to DR
array[178+19] = 26'b00000_01111_000_000_0000000000;//RES-
array[178+20] = 26'b00000_10011_000_000_0000000000;//RES to DR
array[178+21] = 26'b00000_10100_000_000_0000000000;//-DR to RES
array[178+22] = 26'b00000_10011_000_000_0000000000;//RES to DR

array[178+23] = 26'b10111_00000_000_000_0000000000;//DR to TR

array[178+24] = 26'b00001_00101_000_000_0000000000;//PC to AR, PC+TWO
array[178+25] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[178+26] = 26'b00000_01100_000_000_0000000000;//loadOP
array[178+27] = 26'b00000_01001_000_000_0000000000;//OP<<TWO
array[178+28] = 26'b10001_00000_000_000_0000000000;//SP to DR
array[178+29] = 26'b00000_00011_000_000_0000000000;//RES+
array[178+30] = 26'b00000_10011_000_000_0000000000;//RES to DR
array[178+31] = 26'b10010_00000_000_000_0000000000;//DR to SP

array[178+32] = 26'b00000_01110_000_000_0000000000;//SR to OP
array[178+33] = 26'b11000_00100_000_000_0000000000;//SP to AR, incSP
array[178+34] = 26'b00000_10000_000_000_0000000000;//OP to RESULT
array[178+35] = 26'b00101_00000_000_000_0000000000;//RES to mem

array[178+36] = 26'b00000_10001_000_000_0000000000;//SP_STAR to SR

array[178+37] = 26'b01001_00000_000_000_0000000000;//LV to DR
array[178+38] = 26'b11000_00100_000_000_0000000000;//SP to AR, incSP
array[178+39] = 26'b00110_00000_000_000_0000000000;//DR to mem

array[178+40] = 26'b10100_00000_110_000_0000000000;//TR to LV

//return = 218
array[3+215+3] = 26'b00011_00010_000_000_0000000000;//SP_STAR to AR, decSP
array[3+215+4] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[3+215+5] = 26'b00000_01100_000_000_0000000000;//loadOP
array[3+215+6] = 26'b00011_00010_000_000_0000000000;//SP_STAR to AR, decSP
array[3+215+7] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[3+215+8] = 26'b00111_00000_000_000_0000000000;//loadTR
array[3+215+9] = 26'b00011_00010_000_000_0000000000;//SP_STAR to AR, decSP
array[3+215+10] = 26'b00010_00000_000_000_0000000000;//READ MEM;
array[3+215+11] = 26'b00000_11111_000_000_0000000000;//reloadPC from mem

array[3+215+12] = 26'b01001_00000_000_000_0000000000;//LV to DR
array[3+215+13] = 26'b10010_00000_000_000_0000000000;//DR to SP
array[3+215+14] = 26'b10100_00000_000_000_0000000000;//TR to LV


array[3+215+15] = 26'b11000_00100_000_000_0000000000;//SP to AR, incSP
array[3+215+16] = 26'b00000_10000_000_000_0000000000;//OP to RESULT
array[3+215+17] = 26'b00101_00000_110_000_0000000000;//RES to mem


end

assign data=array[address];
endmodule